
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package DORN_Package is

    ----------------------------------------------------------------------------------
    -- Clocks period constants
    ----------------------------------------------------------------------------------

    constant C_UART_PERIOD_NS    : integer range 0 to 200   := 10; -- UART_CLOCK frequency from WFG at 100 MHz
    constant C_UART_BAUDRATE_KBD : integer range 0 to 10000 := 1000; -- Bauderate in [kBit/s], here 1 MBit/s
    constant C_BAUD_CNT_OFFSET   : integer range -15 to 15  := -7; -- Adapt to NX_OSC, can be board dependent
    constant C_PARITY_POL_EVEN   : std_logic                := '0'; -- Even polarity

    constant C_SYSTEM_PERIOD_NS : integer range 0 to 200    := 40; -- MAIN_CLOCK frequency from WFG at 25 MHz, [nanosecond]
    constant C_SYSTEM_PERIOD_PS : integer range 0 to 200000 := C_SYSTEM_PERIOD_NS * 1000; -- [picosecond]

    -- ----------------------------------------------------------------------------------
    -- -- Telecommands (TC) IDs
    -- ----------------------------------------------------------------------------------

    -- constant C_DORN_APID : std_logic_vector(10 downto 0) := 11X"067"; -- DORN_FUSIO_RT Identifier
    -- constant C_UART_EOT  : std_logic_vector(7 downto 0)  := X"55"; -- End Of Transmission

    -- constant C_TC_GET_STATUS   : std_logic_vector(7 downto 0) := X"57";
    -- constant C_TC_START_SC_ACQ : std_logic_vector(7 downto 0) := X"AC";
    -- constant C_TC_PAUSE_SC_ACQ : std_logic_vector(7 downto 0) := X"37";
    -- constant C_TC_RESET_SC_ACQ : std_logic_vector(7 downto 0) := X"B0";
    -- constant C_TC_POWER_OFF    : std_logic_vector(7 downto 0) := X"18";

    -- constant C_TC_LOAD_CONFIG : std_logic_vector(7 downto 0) := X"1C";
    -- constant C_TC_SAVE_CONFIG : std_logic_vector(7 downto 0) := X"5C";

    -- constant C_TC_READ_REGISTER  : std_logic_vector(7 downto 0) := X"D1";
    -- constant C_TC_WRITE_REGISTER : std_logic_vector(7 downto 0) := X"D2";

    -- constant C_TC_FLASH_DUMP  : std_logic_vector(7 downto 0) := X"64";
    -- constant C_TC_FLASH_ERASE : std_logic_vector(7 downto 0) := X"C3";
    -- constant C_TC_FLASH_WRITE : std_logic_vector(7 downto 0) := X"C4";

    -- constant C_TC_EXEC_STATUS_SUCCESS            : std_logic_vector(7 downto 0) := X"22";
    -- constant C_TC_EXEC_STATUS_BAD_APID           : std_logic_vector(7 downto 0) := X"23";
    -- constant C_TC_EXEC_STATUS_BAD_SEQ_FLAGS      : std_logic_vector(7 downto 0) := X"24";
    -- constant C_TC_EXEC_STATUS_BAD_PAYLOAD_LENGTH : std_logic_vector(7 downto 0) := X"25";
    -- constant C_TC_EXEC_STATUS_BAD_EOT            : std_logic_vector(7 downto 0) := X"26";
    -- constant C_TC_EXEC_STATUS_BAD_PCKT_ID        : std_logic_vector(7 downto 0) := X"27";

    -- ----------------------------------------------------------------------------------
    -- -- Telemetries (TM) IDs
    -- ----------------------------------------------------------------------------------

    -- constant C_UART_ERROR   : std_logic_vector(7 downto 0) := X"EE";
    -- constant C_TM_BAD_CMD   : std_logic_vector(7 downto 0) := X"66";
    -- constant C_TM_ACK       : std_logic_vector(7 downto 0) := X"44";
    -- constant C_TM_STATUS    : std_logic_vector(7 downto 0) := X"88";
    -- constant C_TM_DUMP_PCKT : std_logic_vector(7 downto 0) := X"77";

    ----------------------------------------------------------------------------------
    -- TC-TM Flags and Status
    ----------------------------------------------------------------------------------

    type TC_Flags_type is record
        BAD_COMMAND    : std_logic;
        GET_STATUS     : std_logic;
        START_SC_ACQ   : std_logic;
        PAUSE_SC_ACQ   : std_logic;
        RESET_SC_ACQ   : std_logic;
        POWER_OFF      : std_logic;
        LOAD_CONFIG    : std_logic;
        SAVE_CONFIG    : std_logic;
        READ_REGISTER  : std_logic;
        WRITE_REGISTER : std_logic;
        FLASH_DUMP     : std_logic;
        FLASH_ERASE    : std_logic;
        FLASH_WRITE    : std_logic;
    end record TC_Flags_type;

    type TM_Flags_type is record
        ACK_BAD_CMD : std_logic;
        SEND_ACK_OK : std_logic;
        SEND_STATUS : std_logic;
        SEND_DUMP   : std_logic;
    end record TM_Flags_type;

    type HV_Heater_Config_type is record
        COMMAND  : std_logic_vector(11 downto 0); -- DAC Command, calculated by PI control or manual by the user
        MODE     : std_logic_vector(3 downto 0);  -- MSB = 0: On, 1: Off, LSB = 0: Average, 1: HTR_1, 2: HTR_2, 3: Manual
        PI_GAINS : std_logic_vector(7 downto 0);  -- PI Feedback Control, KI & KP
        SETPOINT : std_logic_vector(11 downto 0); -- Heater setpoint, calculated by the user with the transfer function
        MAX_CMD  : std_logic_vector(11 downto 0); -- Heater setpoint, calculated by the user with the transfer function
    end record HV_Heater_Config_type;

    type HV_Commands_Array_type is array (0 to 3) of std_logic_vector(11 downto 0); -- Array 4 x 12

    type TM_Status_type is record
        VERSION       : std_logic_vector(7 downto 0); -- Version number of the bitstream.nxb [0..255]
        MODE          : std_logic_vector(3 downto 0); -- Power-Up (x00), Configuration (x01), Science_Acq (x02), Power-Off(x03)
        HEATER_CFG    : HV_Heater_Config_type;    -- Record (Command, PI_Gains, Setpoint, Mode)
        HV_COMMANDS   : HV_Commands_Array_type;   -- Array 4 x 12: HV_V_A, B, C, D
        HV_FE_On_Off  : std_logic_vector(7 downto 0); -- 4 FE On_Off + 4 HV On_Off
        FPGA_ENABLES  : std_logic_vector(7 downto 0); -- DU_ADC_Meas, Spare, SDRAM, HV, HK, EP, Auto-start_SC, FLASH_Recov
        TEST_PATTERNS : std_logic_vector(3 downto 0); -- 0: No test pattern, 1: Raw and Spectra, 2: P12_Maps, 3: DU_ADC Measures
        DEBUG_PIN_SEL : std_logic_vector(3 downto 0); -- 16 Modes on Debug pins
        DU_ADC_SEL    : std_logic_vector(3 downto 0); -- 12 configurations for displaying DU_ADC data
        STREAM_SEL    : std_logic_vector(3 downto 0); -- 1 Enable and 8 configurations for serial streaming DU_ADC data
    end record TM_Status_type;

    ----------------------------------------------------------------------------------
    -- DORN Registers, max 256 registers, 16 slices of 16 addresses of 16 bits
    -- 8 Slices are used: 0, 1, 2, 3 (Parameters) and C, D, E, F (Measures)
    ----------------------------------------------------------------------------------

    type DORN_Register_Slice_type is array (0 to 15) of std_logic_vector(15 downto 0); -- Array 16 x 16

    -- HV DAC, Power On-Off and Heater Feedback addresses
    constant C_START_REG_HEATER_HV_FE : std_logic_vector(3 downto 0) := X"0"; -- 16 addresses (all used)

    constant C_HEATER_COMMAND_adr    : integer range 0 to 15 := 0;
    constant C_HEATER_MODE_GAINS_adr : integer range 0 to 15 := 1;
    constant C_HEATER_SETPOINT_adr   : integer range 0 to 15 := 2;
    constant C_HEATER_CMD_MAX_adr    : integer range 0 to 15 := 3;
    constant C_FE_2V5_ON_OFF_adr     : integer range 0 to 15 := 4;
    constant C_FE_3V3_ON_OFF_adr     : integer range 0 to 15 := 5; -- C_FE_ON_P7V_DP_adr
    constant C_FE_VCC_7V_ON_OFF_adr  : integer range 0 to 15 := 6; -- C_FE_ON_P7V_M7V_DP10P_adr
    constant C_FE_VSS_7V_ON_OFF_adr  : integer range 0 to 15 := 7; -- C_FE_ON_P7V_M7V_DP20P_adr
    constant C_HV_V_A_COMMAND_adr    : integer range 0 to 15 := 8;
    constant C_HV_V_B_COMMAND_adr    : integer range 0 to 15 := 9;
    constant C_HV_V_C_COMMAND_adr    : integer range 0 to 15 := 10;
    constant C_HV_V_D_COMMAND_adr    : integer range 0 to 15 := 11;
    constant C_HV_A_ON_OFF_adr       : integer range 0 to 15 := 12;
    constant C_HV_B_ON_OFF_adr       : integer range 0 to 15 := 13;
    constant C_HV_C_ON_OFF_adr       : integer range 0 to 15 := 14;
    constant C_HV_D_ON_OFF_adr       : integer range 0 to 15 := 15;

    -- FPGA Configuration addresses
    constant C_START_FPGA_ENABLES : std_logic_vector(3 downto 0) := X"1"; -- 16 addresses (14 used, 2 spare)

    constant C_En_FLASH_Recov_adr    : integer range 0 to 15 := 0;
    constant C_En_AutoStart_SC_adr   : integer range 0 to 15 := 1;
    constant C_En_EP_Generator_adr   : integer range 0 to 15 := 2;
    constant C_En_HK_Generator_adr   : integer range 0 to 15 := 3;
    constant C_En_HV_Generator_adr   : integer range 0 to 15 := 4;
    constant C_Disable_SDRAM_adr     : integer range 0 to 15 := 5;
    constant C_En_Debug_TM_adr       : integer range 0 to 15 := 6;
    constant C_En_DU_ADC_Meas_adr    : integer range 0 to 15 := 7;
    constant C_Test_Patterns_adr     : integer range 0 to 15 := 8;
    constant C_Debug_Pins_Select_adr : integer range 0 to 15 := 9;
    constant C_DU_ADC_Select_adr     : integer range 0 to 15 := 10;
    constant C_Stream_Select_adr     : integer range 0 to 15 := 11;
    constant C_TM_Dead_Time_MSB_adr  : integer range 0 to 15 := 12;
    constant C_TM_Dead_Time_LSB_adr  : integer range 0 to 15 := 13;
    constant C_Spare_5_adr           : integer range 0 to 15 := 14;
    constant C_Spare_6_adr           : integer range 0 to 15 := 15;

    -- DU Configuration addresses
    constant C_START_REG_DU_LDD  : std_logic_vector(3 downto 0) := X"2"; -- 16 addresses (all used)
    constant C_START_REG_DU_THLD : std_logic_vector(3 downto 0) := X"3"; -- 16 addresses (all used)

    ----------------------------------------------------------------------------------
    constant C_END_REG_CONFIG : unsigned(7 downto 0) := X"7F"; -- 128 first addresses
    ----------------------------------------------------------------------------------

    -- FLASH DU_ADC counters
    constant C_START_REG_FLASH_DU_ADC : std_logic_vector(3 downto 0) := X"C"; -- 16 addresses (4 used, 10 spare)

    constant C_FLASH_DUx_ADC_Front_adr : integer range 0 to 15 := 0; -- Area #8
    constant C_FLASH_DUx_ADC_Back_adr  : integer range 0 to 15 := 1; -- Area #9
    constant C_FLASH_DUy_ADC_Front_adr : integer range 0 to 15 := 2; -- Area #10
    constant C_FLASH_DUy_ADC_Back_adr  : integer range 0 to 15 := 3; -- Area #11

    -- FLASH Packets counters
    constant C_START_REG_FLASH_PACKETS : std_logic_vector(3 downto 0) := X"D"; -- 16 addresses (all used)

    constant C_FLASH_PACKETS_Raw_1H_adr  : integer range 0 to 15 := 0; -- Area #0
    constant C_FLASH_PACKETS_Spectra_adr : integer range 0 to 15 := 2; -- Area #1
    constant C_FLASH_PACKETS_P12_Map_adr : integer range 0 to 15 := 4; -- Area #2
    constant C_FLASH_PACKETS_HK_adr      : integer range 0 to 15 := 6; -- Area #3

    constant C_FLASH_PACKETS_Alpha_1H_adr : integer range 0 to 15 := 8; -- Area #4
    constant C_FLASH_PACKETS_Alpha_1L_adr : integer range 0 to 15 := 10; -- Area #5
    constant C_FLASH_PACKETS_Alpha_2_adr  : integer range 0 to 15 := 12; -- Area #6
    constant C_FLASH_PACKETS_Proton12_adr : integer range 0 to 15 := 14; -- Area #7

    -- HK ADC addresses
    constant C_START_REG_HK_VALUES_PART_1 : std_logic_vector(3 downto 0) := X"E"; -- 16 addresses (all used)
    constant C_START_REG_HK_VALUES_PART_2 : std_logic_vector(3 downto 0) := X"F"; -- 16 addresses (all used)

    -- Make sure HK_ID_Temp_Heater_2 < HK_ID_Temp_Heater_1 for sequencing
    constant C_HK_ID_TEMP_HEATER_1 : unsigned(7 downto 0) := X"16"; -- HK_22 = CS2.6
    constant C_HK_ID_TEMP_HEATER_2 : unsigned(7 downto 0) := X"15"; -- HK_21 = CS2.5

    ----------------------------------------------------------------------------------
    -- RIMC SDRAM
    ----------------------------------------------------------------------------------

    -- P12_Map:
    -- Address Part_1 from 0x00_0000 to 0x3F_FFFF  ;  2^22 = 4 194 304 addresses
    -- Address Part_2 from 0x40_0000 to 0x7F_FFFF  ;  2^22 = 4 194 304 addresses
    -- Spectra:
    -- Address Part_1 from 0x80_0000 to 0x83_FFFF  ;  2^18 =   262 144 addresses
    -- Address Part_2 from 0x84_0000 to 0x87_FFFF  ;  2^18 =   262 144 addresses

    -- constant C_SDRAM_END_ADR_ERASING_ALL : unsigned(23 downto 0) := X"87_FE00"; -- 8.9 Mbits to erase

    -- -- 256 beats per burst
    -- constant C_SDRAM_NBR_BEATS_PER_BURST : unsigned(7 downto 0) := X"FF";

    -- -- 16 bursts per packet to make sure the EP_FIFO is never full
    -- constant C_SDRAM_NBR_BURSTS_PER_PACKET : unsigned(3 downto 0) := X"F"; -- 16 bursts of 256 beats of two addresses = 8192 = X"2000" address increment per packet

    -- -- Nbr_Adr / Nbr_Beats / 2 = 2^22 / 2^8 / 2 = 2^13 = 8192 bursts => 512 packets of 16 bursts
    -- constant C_SDRAM_NBR_PACKETS_P12_MAP : unsigned(8 downto 0) := 9X"1FF";
    -- -- Nbr_Adr / Nbr_Beats / 2 = 2^18 / 2^8 / 2 = 2^19  = 512 bursts =>  32 packets of 16 bursts
    -- constant C_SDRAM_NBR_PACKETS_SPECTRA : unsigned(8 downto 0) := 9X"01F";

    ----------------------------------------------------------------------------------
    -- RIMC NAND FLASH
    ----------------------------------------------------------------------------------

    -- -- FLASH Area start addresses, total 4096 blocks
    -- constant C_START_BLOCK_Raw_1H  : std_logic_vector(2 downto 0) := "000"; --  512 blocks, starts at 0x000, ends at 0x1FF
    -- constant C_START_BLOCK_Spectra : std_logic_vector(2 downto 0) := "001"; --  512 blocks, starts at 0x200, ends at 0x3FF
    -- constant C_START_BLOCK_P12_Map : std_logic_vector(1 downto 0) := "01"; --  1024 blocks, starts at 0x400, ends at 0x7FF
    -- constant C_START_BLOCK_HK      : std_logic_vector(3 downto 0) := X"8"; --   256 blocks, starts at 0x800, ends at 0x8FF

    -- constant C_START_BLOCK_Alpha_1H : std_logic_vector(3 downto 0) := X"9"; --  256 blocks, starts at 0x900, ends at 0x9FF
    -- constant C_START_BLOCK_Alpha_1L : std_logic_vector(3 downto 0) := X"A"; --  256 blocks, starts at 0xA00, ends at 0xAFF
    -- constant C_START_BLOCK_Alpha_2  : std_logic_vector(3 downto 0) := X"B"; --  256 blocks, starts at 0xB00, ends at 0xBFF
    -- constant C_START_BLOCK_Proton12 : std_logic_vector(3 downto 0) := X"C"; --  256 blocks, starts at 0xC00, ends at 0xCFF

    -- constant C_START_BLOCK_DUx_ADC_Front : std_logic_vector(4 downto 0) := X"D" & '0'; --  128 blocks, starts at 0xD00, ends at 0xD7F
    -- constant C_START_BLOCK_DUx_ADC_Back  : std_logic_vector(4 downto 0) := X"D" & '1'; --  128 blocks, starts at 0xD80, ends at 0xDFF
    -- constant C_START_BLOCK_DUy_ADC_Front : std_logic_vector(4 downto 0) := X"E" & '0'; --  128 blocks, starts at 0xE00, ends at 0xE7F
    -- constant C_START_BLOCK_DUy_ADC_Back  : std_logic_vector(4 downto 0) := X"E" & '1'; --  128 blocks, starts at 0xE80, ends at 0xEFF

    -- constant C_START_BLOCK_CONFIG : std_logic_vector(7 downto 0) := X"FF"; -- 16 blocks, starts at 0xFF0, ends at 0xFFF

    -- FLASH settings for AXI Stream
    type FLASH_Settings_type is record
        CTYPE  : std_logic_vector(1 downto 0);    -- "00": Erase command, "01": Write command, "10": Read command, "11": Invalid
        BLK    : std_logic_vector(11 downto 0);   -- 4096 blocks in the NAND FLASH module
        PAGE   : std_logic_vector(6 downto 0);    -- 128 pages per block
        CA     : std_logic_vector(12 downto 0);   -- 4096 + 224 = 4320 column addresses per page
        NBDATA : std_logic_vector(23 downto 0);   -- Up to 2^24 - 1 beats of 24-bit data per AXI transaction
    end record FLASH_Settings_type;

    -- -- FLASH data frame tags
    -- constant C_FLASH_START_TAG : std_logic_vector(7 downto 0) := X"AA";
    -- constant C_FLASH_STOP_TAG  : std_logic_vector(7 downto 0) := X"55";

    -- -- FLASH DUMP
    -- constant C_NBR_RAW_SAMPLES   : unsigned(4 downto 0)    := 5D"20"; -- 20 Raw Samples per pulse
    -- constant C_FLASH_DUMP_Size   : integer range 1 to 11   := 10; -- Output FIFO DUMP size
    -- constant C_FLASH_DUMP_Packet : integer range 1 to 2047 := 2 ** C_FLASH_DUMP_Size - 1; -- 1024 data of 24 bits per dump packet maximum
    -- constant C_FIFO_EVENTS_Size  : integer range 1 to 11   := C_FLASH_DUMP_Size + 1; -- 2048 data per FIFO maximum before saturation

    -- -- 1024 data are written per dump packet in a page
    -- constant C_FLASH_NBDATA_Pckt : std_logic_vector(23 downto 0) := std_logic_vector(to_unsigned(C_FLASH_DUMP_Packet, 24)); -- NBDATA = 0x00_03FF
    -- -- 128 first registers addresses data are written in the FLASH
    -- constant C_NBDATA_CONFIG     : std_logic_vector(23 downto 0) := std_logic_vector(resize(C_END_REG_CONFIG, 24));
    ----------------------------------------------------------------------------------
    -- Event Processor
    ----------------------------------------------------------------------------------


	
    type Array_8x6_type is array (0 to 7) of std_logic_vector(5 downto 0); -- Array 8 x 6
    type Array_8x16_type is array (0 to 7) of std_logic_vector(15 downto 0); -- Array 8 x 16
	
	type Array_4x31_type is array (0 to 3) of signed(31 downto 0); -- Array 8 x 16
	type Array_8x31_type is array (0 to 7) of signed(31 downto 0); -- Array 8 x 16
	
	type Array_4x16_type is array (0 to 3) of std_logic_vector(15 downto 0); -- Array 4 x 16
	
    -- constant C_DU_ADC_LLD_DEFAULT  : std_logic_vector(15 downto 0) := X"7777"; -- DEBUG value
    -- constant C_DU_THLD_1H_DEFAULT  : std_logic_vector(15 downto 0) := X"8888"; -- DEBUG value
    -- constant C_DU_THLD_RAW_DEFAULT : std_logic_vector(15 downto 0) := X"9999"; -- DEBUG value

    -- EP_Data Structure for Events:
    -- # Bit  # Size    # Name          # Description
    -- 23:       1       Time_Flag       0: Energy value, standard header
    -- 22:       1       Raw_Flag        0: Events, 1: Raw Samples
    -- 21..20    2       Event_Type      "00": Alpha_1H, "01": Alpha_1L, "10": Alpha_2, "11": Proton12
    -- 19..16    4       ADC_ID          16 Detectors ADC ID, 2 per DU, Even = Front, Odd = Back
    -- 15..0:   16       Energy Value    16-bit signed value

    -- EP_Data Structure for Timestamp:
    -- # Bit  # Size    # Name          # Description
    -- 23:       1       Time_Flag       1: Timestamp, no header
    -- 22..0:   23       Time Value      23-bit unsigned value, 1 LSB = 1 �s, max ~8.39s

    ----------------------------------------------------------------------------------
    -- Front-end Power, HV_DAC, HK_ADC, DU_TEMP_ADC, Heater Feedback
    ----------------------------------------------------------------------------------

    -- HV_1 max voltage = -110V <=> 3.3V    DAC => HV_1 Command = -70V <=> V_Command = 70 / 110 * 3.3 = 2.10V
    -- HV_2 max voltage =  -66V <=> 3.3V    DAC => HV_2 Command = -20V <=> V_Command = 20 /  66 * 3.3 = 1.00V

    -- DAC Full scale : X"FFF" => 3.2992 V
    -- Vout = N_Command * 3.3V / 4096
    -- N_HV1_CMD = round_up(2.10 * 4096 / 3.3) = X"0A2F"
    -- N_HV1_CMD = round_up(1.00 * 4096 / 3.3) = X"04DA"

    -- constant C_HV_HEATER_COMMAND_MAX : std_logic_vector(11 downto 0) := X"FFF"; -- 3.2992 V <=> 88.0�C
    -- constant C_HV_HEATER_PI_KI       : std_logic_vector(3 downto 0)  := X"2"; -- => Ki = 2^(-2) = 1/4
    -- constant C_HV_HEATER_PI_KP       : std_logic_vector(3 downto 0)  := X"4"; -- => Kp = 4 V/V

    ----------------------------------------------------------------------------------
    -- Memory Init Data
    ----------------------------------------------------------------------------------

    --    constant C_RAM_Init_2kx24 : string := ( -- All zeros
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000," &
    --"000000000000000000000000,000000000000000000000000,000000000000000000000000,000000000000000000000000");

    --    constant C_RBF_Init : string := (   -- All zeros
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000," &
    --    "0000000000000000,0000000000000000," & "0000000000000000,0000000000000000");

end package DORN_Package;
