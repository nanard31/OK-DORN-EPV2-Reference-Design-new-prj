Library ieee;
use ieee.std_logic_1164.all;

entity Coeff_Table is
	port(address : in  integer range 0 to 255;
		 data    : out integer range 0 to 131071
	);
end entity Coeff_Table;

architecture behavioral of Coeff_Table is
	type Table is array (0 to 255) of integer range 0 to 131071;
	constant Table_Value : Table := (
 65602 ,
 65607 ,
 65613 ,
 65619 ,
 65625 ,
 65631 ,
 65637 ,
 65643 ,
 65649 ,
 65655 ,
 65661 ,
 65668 ,
 65676 ,
 65683 ,
 65691 ,
 65699 ,
 65707 ,
 65715 ,
 65723 ,
 65732 ,
 65740 ,
 65749 ,
 65758 ,
 65767 ,
 65777 ,
 65787 ,
 65797 ,
 65808 ,
 65819 ,
 65830 ,
 65841 ,
 65852 ,
 65863 ,
 65874 ,
 65885 ,
 65896 ,
 65908 ,
 65919 ,
 65931 ,
 65943 ,
 65956 ,
 65968 ,
 65981 ,
 65994 ,
 66008 ,
 66021 ,
 66035 ,
 66049 ,
 66063 ,
 66077 ,
 66091 ,
 66105 ,
 66119 ,
 66133 ,
 66147 ,
 66160 ,
 66173 ,
 66186 ,
 66199 ,
 66211 ,
 66223 ,
 66234 ,
 66245 ,
 66255 ,
 66265 ,
 66274 ,
 66282 ,
 66289 ,
 66296 ,
 66302 ,
 66307 ,
 66311 ,
 66314 ,
 66317 ,
 66318 ,
 66318 ,
 66317 ,
 66314 ,
 66311 ,
 66306 ,
 66300 ,
 66293 ,
 66284 ,
 66274 ,
 66262 ,
 66249 ,
 66234 ,
 66218 ,
 66199 ,
 66180 ,
 66158 ,
 66135 ,
 66110 ,
 66083 ,
 66054 ,
 66023 ,
 65990 ,
 65955 ,
 65918 ,
 65879 ,
 65838 ,
 65794 ,
 65748 ,
 65700 ,
 65649 ,
 65597 ,
 65541 ,
 65483 ,
 65423 ,
 65360 ,
 65294 ,
 65226 ,
 65155 ,
 65081 ,
 65005 ,
 64926 ,
 64843 ,
 64758 ,
 64670 ,
 64579 ,
 64485 ,
 64388 ,
 64287 ,
 64183 ,
 64077 ,
 63966 ,
 63853 ,
 63736 ,
 68903 ,
 68779 ,
 68658 ,
 68542 ,
 68429 ,
 68321 ,
 68216 ,
 68114 ,
 68016 ,
 67922 ,
 67830 ,
 67743 ,
 67658 ,
 67576 ,
 67498 ,
 67422 ,
 67349 ,
 67280 ,
 67212 ,
 67148 ,
 67086 ,
 67026 ,
 66969 ,
 66914 ,
 66861 ,
 66810 ,
 66762 ,
 66715 ,
 66670 ,
 66628 ,
 66586 ,
 66547 ,
 66509 ,
 66472 ,
 66437 ,
 66403 ,
 66370 ,
 66339 ,
 66308 ,
 66279 ,
 66250 ,
 66223 ,
 66196 ,
 66169 ,
 66143 ,
 66118 ,
 66093 ,
 66069 ,
 66044 ,
 66020 ,
 65996 ,
 65972 ,
 65947 ,
 65923 ,
 65898 ,
 65873 ,
 65848 ,
 65822 ,
 65797 ,
 65774 ,
 65752 ,
 65732 ,
 65716 ,
 65703 ,
 65692 ,
 65682 ,
 65674 ,
 65667 ,
 65659 ,
 65651 ,
 65644 ,
 65637 ,
 65630 ,
 65623 ,
 65617 ,
 65611 ,
 65605 ,
 65599 ,
 65594 ,
 65590 ,
 65585 ,
 65581 ,
 65577 ,
 65574 ,
 65570 ,
 65566 ,
 65563 ,
 65559 ,
 65556 ,
 65553 ,
 65550 ,
 65547 ,
 65545 ,
 65543 ,
 65541 ,
 65540 ,
 65539 ,
 65539 ,
 65538 ,
 65538 ,
 65537 ,
 65536 ,
 65536 ,
 65535 ,
 65535 ,
 65535 ,
 65536 ,
 65537 ,
 65539 ,
 65541 ,
 65543 ,
 65545 ,
 65547 ,
 65548 ,
 65550 ,
 65553 ,
 65555 ,
 65557 ,
 65560 ,
 65564 ,
 65567 ,
 65571 ,
 65575 ,
 65579 ,
 65583 ,
 65587 ,
 65592 ,
 65597 
); -- bit 17 is 0 or 1 decimal bit 16 to 0 are mantis 2^negative

begin

data <= Table_Value(address);
end architecture behavioral;
--C:\Projets\DORN\Pulse_Processor\OpalKelly\OK-DORN-RAW-PeakAndHold\DDR3Loader\DDR3Loader.runs\impl_1

--65888,
--65862,
--65838,
--65815,
--65793,
--65772,
--65751,
--65732,
--65714,
--65696,
--65680,
--65664,
--65650,
--65636,
--65623,
--65611,
--65601,
--65591,
--65581,
--65573,
--65566,
--65560,
--65554,
--65549,
--65546,
--65543,
--65541,
--65540,
--65539,
--65540,
--65541,
--65544,
--65547,
--65550,
--65555,
--65561,
--65567,
--65574,
--65582,
--65591,
--65601,
--65611,
--65623,
--65635,
--65648,
--65661,
--65676,
--65691,
--65707,
--65724,
--65741,
--65759,
--65778,
--65798,
--65819,
--65840,
--65862,
--65885,
--65909,
--65933